module auth_login

enum AuthProvider {
	google
	github
	// Adicione outros provedores de autenticação aqui
}
